library verilog;
use verilog.vl_types.all;
entity LPM_MEMORY_INITIALIZATION is
end LPM_MEMORY_INITIALIZATION;
