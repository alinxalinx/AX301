library verilog;
use verilog.vl_types.all;
entity shift_tb is
end shift_tb;
