library verilog;
use verilog.vl_types.all;
entity led_test_tb is
end led_test_tb;
